/*  This file is part of JTS16.
    JTS16 program is free software: you can redistribute it and/or modify
    it under the terms of the GNU General Public License as published by
    the Free Software Foundation, either version 3 of the License, or
    (at your option) any later version.

    JTS16 program is distributed in the hope that it will be useful,
    but WITHOUT ANY WARRANTY; without even the implied warranty of
    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
    GNU General Public License for more details.

    You should have received a copy of the GNU General Public License
    along with JTS16.  If not, see <http://www.gnu.org/licenses/>.

    Author: Jose Tejada Gomez. Twitter: @topapate
    Version: 1.0
    Date: 5-7-2021 */

`ifndef NOSOUND

module jts16b_snd(
    input                rst,
    input                clk,

    input                cen_snd,   // 5MHz -- jumper to select 5 or 4MHz
    input                cen_fm,    // 4MHz
    input                cen_fm2,   // 2MHz
    input                cen_pcm,   // 0.640

    input                sound_en,
    // options
    input         [ 1:0] fxlevel,
    input                enable_fm,
    input                enable_psg,

    input         [ 7:0] latch,
    output               ack,

    // Mapper device 315-5195
    output               mapper_rd,
    output               mapper_wr,
    output [7:0]         mapper_din,
    input  [7:0]         mapper_dout,
    input                mapper_obf, // pbf signal == buffer full ?

    // ROM
    output    reg [18:0] rom_addr,
    output    reg        rom_cs,
    input         [ 7:0] rom_data,
    input                rom_ok,

    // Sound output
    output signed [15:0] snd,
    output               sample,
    output               peak
);

localparam [7:0] FMGAIN=8'h10;

wire [15:0] A;
reg         fm_cs, mapper_cs, ram_cs, bank_cs;
wire        mreq_n, iorq_n, int_n;
wire        WRn;
reg  [ 7:0] din, pcm_cmd, pcmgain;
reg         rom_ok2;
wire        rom_good, cmd_cs;
wire [ 7:0] dout, fm_dout, ram_dout;
wire        nmi_n, pcm_busyn,
            wr_n, rd_n;
reg         pcm_mdn, pcm_rst;
reg  [ 5:0] rom_msb;


wire signed [15:0] fm_left, fm_right, mixed;
wire signed [ 8:0] pcm_raw, pcm_snd;
wire [7:0] fmgain;

assign snd = sound_en ? mixed : 16'd0;

assign rom_good = rom_ok2 & rom_ok;
assign ack      = mapper_cs;
assign cmd_cs   = !iorq_n && A[7:6]==2 && !wr_n; // 80
assign fmgain   = enable_fm ? FMGAIN : 0;

assign mapper_rd   = mapper_cs && !rd_n;
assign mapper_wr   = mapper_cs && !wr_n;
assign mapper_dout = cpu_dout;

// ROM bank address
always @(*) begin
    rom_addr = { 6'd0, A[14:0] };
    if( bank_cs ) begin
        // For board type 171-5358
        rom_addr[15:14] = rom_msb[1:0];
        casez( rom_msb[5:2] ) // A11-A8 refer to the ROM label in the PCB:
            4'b1???: rom_addr[17:16] = 3; // A11 at top
            4'b01??: rom_addr[17:16] = 2; // A10
            4'b001?: rom_addr[17:16] = 1; // A9
            4'b0001: rom_addr[17:16] = 0; // A8
        endcase
    end
end

// PCM volume
always @(posedge clk ) begin
    case( fxlevel )
        2'd0: pcmgain <= 8'h04;
        2'd1: pcmgain <= 8'h06;
        2'd2: pcmgain <= 8'h08;
        2'd3: pcmgain <= 8'h0C;
    endcase
    if( !enable_psg ) pcmgain <= 0;
end

always @(*) begin
    bank_cs = !mreq_n && (A[15:12]>=8 && A[15:12]<4'he);
    // Port Map
    if( !iorq_n ) begin
        case( A[7:6] )
            0: fm_cs     = 1;
            1: misc_cs   = 1;
            2: upd_st_cs = 1;
            3: mapper_cs = 1;
        endcase
    end else begin
        mapper_cs = (!mreq_n &&  A[15:12]==4'he && A[11]) // e800
    end
end

always @(posedge clk) begin
    ram_cs   <=  !mreq_n && &A[15:11];
    rom_cs   <=  (!mreq_n && !A[15]) || bank_cs;
    rom_ok2  <= rom_ok;
    if( cmd_cs ) pcm_cmd <= dout;

    din      <= rom_cs    ? rom_data : (
                ram_cs    ? ram_dout : (
                fm_cs     ? fm_dout  : (
                mapper_cs ? mapper_dout : (
                    8'hff ))));
end

always @(posedge clk, posedge rst) begin
    if( rst ) begin
        rom_msb <= 0;
    end else if(misc_cs) begin
        rom_msb <= cpu_dout[5:0];
        pcm_rst <= ~cpu_dout[6];
        pcm_mdn <= cpu_dout[7];
    end
end

jtframe_mixer #(.W2(9)) u_mixer(
    .rst    ( rst       ),
    .clk    ( clk       ),
    .cen    ( 1'b1      ),
    // input signals
    .ch0    ( fm_left   ),
    .ch1    ( fm_right  ),
    .ch2    ( pcm_snd   ),
    .ch3    ( 16'd0     ),
    // gain for each channel in 4.4 fixed point format
    .gain0  ( fmgain    ),
    .gain1  ( fmgain    ),
    .gain2  ( pcmgain   ),
    .gain3  ( 8'h00     ),
    .mixed  ( mixed     ),
    .peak   ( peak      )
);

jtframe_ff u_ff(
    .rst    ( rst       ),
    .clk    ( clk       ),
    .cen    ( 1'b1      ),
    .din    ( 1'b1      ),
    .q      (           ),
    .qn     ( int_n     ),
    .set    ( 1'b0      ),    // active high
    .clr    ( mapper_cs  ),    // active high
    .sigedge( mapper_obf ) // signal whose edge will trigger the FF
);

jtframe_sysz80 #(.RAM_AW(11)) u_cpu(
    .rst_n      ( ~rst        ),
    .clk        ( clk         ),
    .cen        ( cen_snd     ),
    .cpu_cen    (             ),
    .int_n      ( int_n       ),
    .nmi_n      ( nmi_n       ),
    .busrq_n    ( 1'b1        ),
    .m1_n       (             ),
    .mreq_n     ( mreq_n      ),
    .iorq_n     ( iorq_n      ),
    .rd_n       ( rd_n        ),
    .wr_n       ( wr_n        ),
    .rfsh_n     (             ),
    .halt_n     (             ),
    .busak_n    (             ),
    .A          ( A           ),
    .cpu_din    ( din         ),
    .cpu_dout   ( dout        ),
    .ram_dout   ( ram_dout    ),
    // manage access to ROM data from SDRAM
    .ram_cs     ( ram_cs      ),
    .rom_cs     ( rom_cs      ),
    .rom_ok     ( rom_good    )
);

//
//  YM2151 output port
//
//  D1 = /RESET line on 7751
//  D0 = /IRQ line on 7751
//

jt51 u_jt51(
    .rst        ( rst       ), // reset
    .clk        ( clk       ), // main clock
    .cen        ( cen_fm    ),
    .cen_p1     ( cen_fm2   ),
    .cs_n       ( !fm_cs    ), // chip select
    .wr_n       ( wr_n      ), // write
    .a0         ( A[0]      ),
    .din        ( dout      ), // data in
    .dout       ( fm_dout   ), // data out
    .ct1        (           ),
    .ct2        (           ),
    .irq_n      ( int_n     ),  // I do not synchronize this signal
    // Low resolution output (same as real chip)
    .sample     ( sample    ), // marks new output sample
    .left       (           ),
    .right      (           ),
    // Full resolution output
    .xleft      ( fm_left   ),
    .xright     ( fm_right  ),
    // unsigned outputs for sigma delta converters, full resolution
    .dacleft    (           ),
    .dacright   (           )
);

jt7759 u_pcm(
    .rst        ( pcm_rst   ), // reset
    .clk        ( clk       ), // main clock
    .cen        ( cen_pcm   ),  // 640kHz
    .stn        ( 1'b1      ),  // STart (active low)
    .cs         ( pcm_cs    ),
    .mdn        ( pcm_mdn   ),  // MODE: 1 for stand alone mode, 0 for slave mode
    .busyn      ( pcm_busyn ),
    // CPU interface
    .wrn        ( wr_n      ),  // for slave mode only
    .din        ( cpu_dout  ),
    .drq        ( nmi_n     ),
    // ROM interface
    .rom_cs     (           ),      // equivalent to DRQn in original chip
    .rom_addr   (           ),
    .rom_data   (           ),
    .rom_ok     ( 1'b0      ),
    // Sound output
    .sound      ( pcm_raw   )
);

// where a = exp(-wc/T ), a<1
// wc = radian frequency

wire [3:0] pole_a = 4'd10; // pole at 4kHz

jtframe_pole #(.WS(9)) u_pole(
    .rst        ( rst       ),
    .clk        ( clk       ),
    .sample     ( sample    ),      // uses the YM2151 as sampling signal
    .a          ( pole_a    ),
    .sin        ( pcm_raw   ),
    .sout       ( pcm_snd   )
);

endmodule

`endif